module Module;

endmodule
